/* Automatically generated from https://wokwi.com/projects/380408823952452609 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_380408823952452609(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = rst_n;
  wire net3 = ui_in[0];
  wire net4 = ui_in[1];
  wire net5 = ui_in[2];
  wire net6 = ui_in[3];
  wire net7 = ui_in[4];
  wire net8;
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16 = 1'b0;
  wire net17 = 1'b1;
  wire net18 = 1'b1;
  wire net19 = 1'b0;
  wire net20 = 1'b1;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42 = 1'b1;
  wire net43;
  wire net44 = 1'b0;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51 = 1'b0;
  wire net52;
  wire net53 = 1'b1;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60 = 1'b1;
  wire net61 = 1'b0;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69 = 1'b0;
  wire net70 = 1'b1;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78 = 1'b1;
  wire net79 = 1'b0;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87 = 1'b1;
  wire net88 = 1'b0;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96 = 1'b1;
  wire net97 = 1'b0;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105 = 1'b0;
  wire net106 = 1'b1;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114 = 1'b0;
  wire net115 = 1'b1;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123 = 1'b0;
  wire net124 = 1'b1;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132 = 1'b1;
  wire net133 = 1'b0;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141 = 1'b0;
  wire net142;
  wire net143 = 1'b1;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150 = 1'b1;
  wire net151 = 1'b0;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159 = 1'b0;
  wire net160;
  wire net161 = 1'b1;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168 = 1'b1;
  wire net169;
  wire net170;
  wire net171;
  wire net172 = 1'b0;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177 = 1'b1;
  wire net178;
  wire net179 = 1'b0;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186 = 1'b1;
  wire net187;
  wire net188 = 1'b0;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195 = 1'b0;
  wire net196;
  wire net197;
  wire net198 = 1'b1;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204 = 1'b1;
  wire net205 = 1'b0;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213 = 1'b0;
  wire net214;
  wire net215 = 1'b1;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222 = 1'b0;
  wire net223;
  wire net224 = 1'b1;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231 = 1'b0;
  wire net232;
  wire net233 = 1'b1;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240 = 1'b1;
  wire net241 = 1'b0;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249 = 1'b1;
  wire net250 = 1'b0;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258 = 1'b0;
  wire net259 = 1'b1;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267 = 1'b1;
  wire net268;
  wire net269 = 1'b0;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276 = 1'b0;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284 = 1'b0;
  wire net285;
  wire net286 = 1'b1;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293 = 1'b0;
  wire net294;
  wire net295;
  wire net296;
  wire net297 = 1'b1;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302 = 1'b0;
  wire net303;
  wire net304;
  wire net305;
  wire net306 = 1'b1;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311 = 1'b0;
  wire net312 = 1'b1;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320 = 1'b0;
  wire net321 = 1'b1;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;

  assign uo_out[0] = net8;
  assign uo_out[1] = net9;
  assign uo_out[2] = net10;
  assign uo_out[3] = net11;
  assign uo_out[4] = net12;
  assign uo_out[5] = net13;
  assign uo_out[6] = net14;
  assign uo_out[7] = net15;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  dffsr_cell flop1 (
    .d (net21),
    .clk (net1),
    .r (net22),
    .q (net23),
    .notq (net21)
  );
  dffsr_cell flop2 (
    .d (net24),
    .clk (net23),
    .r (net22),
    .q (net25),
    .notq (net24)
  );
  dffsr_cell flop3 (
    .d (net26),
    .clk (net25),
    .r (net22),
    .q (net27),
    .notq (net26)
  );
  not_cell not1 (
    .in (net2),
    .out (net22)
  );
  and_cell and1 (
    .a (net28),
    .b (net29),
    .out (net8)
  );
  and_cell and2 (
    .a (net23),
    .b (net29),
    .out (net9)
  );
  not_cell not2 (
    .in (net23),
    .out (net28)
  );
  and_cell and3 (
    .a (net30),
    .b (net31),
    .out (net10)
  );
  and_cell and4 (
    .a (net23),
    .b (net31),
    .out (net11)
  );
  not_cell not3 (
    .in (net23),
    .out (net30)
  );
  and_cell and5 (
    .a (net32),
    .b (net33),
    .out (net12)
  );
  and_cell and6 (
    .a (net23),
    .b (net33),
    .out (net13)
  );
  not_cell not4 (
    .in (net23),
    .out (net32)
  );
  and_cell and7 (
    .a (net34),
    .b (net35),
    .out (net14)
  );
  and_cell and8 (
    .a (net23),
    .b (net35),
    .out (net15)
  );
  not_cell not5 (
    .in (net23),
    .out (net34)
  );
  and_cell and9 (
    .a (net36),
    .b (net37),
    .out (net29)
  );
  and_cell and10 (
    .a (net25),
    .b (net37),
    .out (net31)
  );
  not_cell not6 (
    .in (net25),
    .out (net36)
  );
  and_cell and11 (
    .a (net38),
    .b (net39),
    .out (net33)
  );
  and_cell and12 (
    .a (net25),
    .b (net39),
    .out (net35)
  );
  not_cell not7 (
    .in (net25),
    .out (net38)
  );
  and_cell and13 (
    .a (net40),
    .b (net41),
    .out (net37)
  );
  and_cell and14 (
    .a (net27),
    .b (net41),
    .out (net39)
  );
  not_cell not8 (
    .in (net27),
    .out (net40)
  );
  mux_cell mux1 (
    .a (net42),
    .b (net42),
    .sel (net23),
    .out (net43)
  );
  mux_cell mux2 (
    .a (net42),
    .b (net44),
    .sel (net23),
    .out (net45)
  );
  mux_cell mux3 (
    .a (net42),
    .b (net42),
    .sel (net23),
    .out (net46)
  );
  mux_cell mux4 (
    .a (net42),
    .b (net44),
    .sel (net23),
    .out (net47)
  );
  mux_cell mux5 (
    .a (net43),
    .b (net45),
    .sel (net25),
    .out (net48)
  );
  mux_cell mux6 (
    .a (net46),
    .b (net47),
    .sel (net25),
    .out (net49)
  );
  mux_cell mux7 (
    .a (net48),
    .b (net49),
    .sel (net27),
    .out (net50)
  );
  mux_cell mux8 (
    .a (net51),
    .b (net51),
    .sel (net23),
    .out (net52)
  );
  mux_cell mux9 (
    .a (net53),
    .b (net53),
    .sel (net23),
    .out (net54)
  );
  mux_cell mux10 (
    .a (net53),
    .b (net53),
    .sel (net23),
    .out (net55)
  );
  mux_cell mux11 (
    .a (net53),
    .b (net51),
    .sel (net23),
    .out (net56)
  );
  mux_cell mux12 (
    .a (net52),
    .b (net54),
    .sel (net25),
    .out (net57)
  );
  mux_cell mux13 (
    .a (net55),
    .b (net56),
    .sel (net25),
    .out (net58)
  );
  mux_cell mux14 (
    .a (net57),
    .b (net58),
    .sel (net27),
    .out (net59)
  );
  mux_cell mux15 (
    .a (net60),
    .b (net61),
    .sel (net23),
    .out (net62)
  );
  mux_cell mux16 (
    .a (net61),
    .b (net60),
    .sel (net23),
    .out (net63)
  );
  mux_cell mux17 (
    .a (net60),
    .b (net60),
    .sel (net23),
    .out (net64)
  );
  mux_cell mux18 (
    .a (net61),
    .b (net61),
    .sel (net23),
    .out (net65)
  );
  mux_cell mux19 (
    .a (net62),
    .b (net63),
    .sel (net25),
    .out (net66)
  );
  mux_cell mux20 (
    .a (net64),
    .b (net65),
    .sel (net25),
    .out (net67)
  );
  mux_cell mux21 (
    .a (net66),
    .b (net67),
    .sel (net27),
    .out (net68)
  );
  mux_cell mux22 (
    .a (net69),
    .b (net70),
    .sel (net23),
    .out (net71)
  );
  mux_cell mux23 (
    .a (net70),
    .b (net70),
    .sel (net23),
    .out (net72)
  );
  mux_cell mux24 (
    .a (net70),
    .b (net69),
    .sel (net23),
    .out (net73)
  );
  mux_cell mux25 (
    .a (net70),
    .b (net69),
    .sel (net23),
    .out (net74)
  );
  mux_cell mux26 (
    .a (net71),
    .b (net72),
    .sel (net25),
    .out (net75)
  );
  mux_cell mux27 (
    .a (net73),
    .b (net74),
    .sel (net25),
    .out (net76)
  );
  mux_cell mux28 (
    .a (net75),
    .b (net76),
    .sel (net27),
    .out (net77)
  );
  mux_cell mux29 (
    .a (net78),
    .b (net79),
    .sel (net23),
    .out (net80)
  );
  mux_cell mux30 (
    .a (net79),
    .b (net78),
    .sel (net23),
    .out (net81)
  );
  mux_cell mux31 (
    .a (net78),
    .b (net78),
    .sel (net23),
    .out (net82)
  );
  mux_cell mux32 (
    .a (net78),
    .b (net79),
    .sel (net23),
    .out (net83)
  );
  mux_cell mux33 (
    .a (net80),
    .b (net81),
    .sel (net25),
    .out (net84)
  );
  mux_cell mux34 (
    .a (net82),
    .b (net83),
    .sel (net25),
    .out (net85)
  );
  mux_cell mux35 (
    .a (net84),
    .b (net85),
    .sel (net27),
    .out (net86)
  );
  mux_cell mux36 (
    .a (net87),
    .b (net88),
    .sel (net23),
    .out (net89)
  );
  mux_cell mux37 (
    .a (net88),
    .b (net88),
    .sel (net23),
    .out (net90)
  );
  mux_cell mux38 (
    .a (net87),
    .b (net87),
    .sel (net23),
    .out (net91)
  );
  mux_cell mux39 (
    .a (net87),
    .b (net88),
    .sel (net23),
    .out (net92)
  );
  mux_cell mux40 (
    .a (net89),
    .b (net90),
    .sel (net25),
    .out (net93)
  );
  mux_cell mux41 (
    .a (net91),
    .b (net92),
    .sel (net25),
    .out (net94)
  );
  mux_cell mux42 (
    .a (net93),
    .b (net94),
    .sel (net27),
    .out (net95)
  );
  mux_cell mux43 (
    .a (net96),
    .b (net97),
    .sel (net23),
    .out (net98)
  );
  mux_cell mux44 (
    .a (net96),
    .b (net96),
    .sel (net23),
    .out (net99)
  );
  mux_cell mux45 (
    .a (net96),
    .b (net96),
    .sel (net23),
    .out (net100)
  );
  mux_cell mux46 (
    .a (net97),
    .b (net97),
    .sel (net23),
    .out (net101)
  );
  mux_cell mux47 (
    .a (net98),
    .b (net99),
    .sel (net25),
    .out (net102)
  );
  mux_cell mux48 (
    .a (net100),
    .b (net101),
    .sel (net25),
    .out (net103)
  );
  mux_cell mux49 (
    .a (net102),
    .b (net103),
    .sel (net27),
    .out (net104)
  );
  mux_cell mux50 (
    .a (net105),
    .b (net106),
    .sel (net23),
    .out (net107)
  );
  mux_cell mux51 (
    .a (net106),
    .b (net105),
    .sel (net23),
    .out (net108)
  );
  mux_cell mux52 (
    .a (net106),
    .b (net106),
    .sel (net23),
    .out (net109)
  );
  mux_cell mux53 (
    .a (net106),
    .b (net105),
    .sel (net23),
    .out (net110)
  );
  mux_cell mux54 (
    .a (net107),
    .b (net108),
    .sel (net25),
    .out (net111)
  );
  mux_cell mux55 (
    .a (net109),
    .b (net110),
    .sel (net25),
    .out (net112)
  );
  mux_cell mux56 (
    .a (net111),
    .b (net112),
    .sel (net27),
    .out (net113)
  );
  mux_cell mux57 (
    .a (net114),
    .b (net115),
    .sel (net23),
    .out (net116)
  );
  mux_cell mux58 (
    .a (net115),
    .b (net114),
    .sel (net23),
    .out (net117)
  );
  mux_cell mux59 (
    .a (net114),
    .b (net114),
    .sel (net23),
    .out (net118)
  );
  mux_cell mux60 (
    .a (net114),
    .b (net114),
    .sel (net23),
    .out (net119)
  );
  mux_cell mux61 (
    .a (net116),
    .b (net117),
    .sel (net25),
    .out (net120)
  );
  mux_cell mux62 (
    .a (net118),
    .b (net119),
    .sel (net25),
    .out (net121)
  );
  mux_cell mux63 (
    .a (net120),
    .b (net121),
    .sel (net27),
    .out (net122)
  );
  mux_cell mux64 (
    .a (net123),
    .b (net124),
    .sel (net23),
    .out (net125)
  );
  mux_cell mux65 (
    .a (net124),
    .b (net124),
    .sel (net23),
    .out (net126)
  );
  mux_cell mux66 (
    .a (net123),
    .b (net123),
    .sel (net23),
    .out (net127)
  );
  mux_cell mux67 (
    .a (net123),
    .b (net123),
    .sel (net23),
    .out (net128)
  );
  mux_cell mux68 (
    .a (net125),
    .b (net126),
    .sel (net25),
    .out (net129)
  );
  mux_cell mux69 (
    .a (net127),
    .b (net128),
    .sel (net25),
    .out (net130)
  );
  mux_cell mux70 (
    .a (net129),
    .b (net130),
    .sel (net27),
    .out (net131)
  );
  mux_cell mux71 (
    .a (net132),
    .b (net133),
    .sel (net23),
    .out (net134)
  );
  mux_cell mux72 (
    .a (net132),
    .b (net133),
    .sel (net23),
    .out (net135)
  );
  mux_cell mux73 (
    .a (net132),
    .b (net132),
    .sel (net23),
    .out (net136)
  );
  mux_cell mux74 (
    .a (net132),
    .b (net133),
    .sel (net23),
    .out (net137)
  );
  mux_cell mux75 (
    .a (net134),
    .b (net135),
    .sel (net25),
    .out (net138)
  );
  mux_cell mux76 (
    .a (net136),
    .b (net137),
    .sel (net25),
    .out (net139)
  );
  mux_cell mux77 (
    .a (net138),
    .b (net139),
    .sel (net27),
    .out (net140)
  );
  mux_cell mux78 (
    .a (net141),
    .b (net141),
    .sel (net23),
    .out (net142)
  );
  mux_cell mux79 (
    .a (net141),
    .b (net143),
    .sel (net23),
    .out (net144)
  );
  mux_cell mux80 (
    .a (net143),
    .b (net143),
    .sel (net23),
    .out (net145)
  );
  mux_cell mux81 (
    .a (net141),
    .b (net141),
    .sel (net23),
    .out (net146)
  );
  mux_cell mux82 (
    .a (net142),
    .b (net144),
    .sel (net25),
    .out (net147)
  );
  mux_cell mux83 (
    .a (net145),
    .b (net146),
    .sel (net25),
    .out (net148)
  );
  mux_cell mux84 (
    .a (net147),
    .b (net148),
    .sel (net27),
    .out (net149)
  );
  mux_cell mux85 (
    .a (net150),
    .b (net151),
    .sel (net23),
    .out (net152)
  );
  mux_cell mux86 (
    .a (net150),
    .b (net151),
    .sel (net23),
    .out (net153)
  );
  mux_cell mux87 (
    .a (net150),
    .b (net151),
    .sel (net23),
    .out (net154)
  );
  mux_cell mux88 (
    .a (net150),
    .b (net151),
    .sel (net23),
    .out (net155)
  );
  mux_cell mux89 (
    .a (net152),
    .b (net153),
    .sel (net25),
    .out (net156)
  );
  mux_cell mux90 (
    .a (net154),
    .b (net155),
    .sel (net25),
    .out (net157)
  );
  mux_cell mux91 (
    .a (net156),
    .b (net157),
    .sel (net27),
    .out (net158)
  );
  mux_cell mux92 (
    .a (net159),
    .b (net159),
    .sel (net23),
    .out (net160)
  );
  mux_cell mux93 (
    .a (net161),
    .b (net159),
    .sel (net23),
    .out (net162)
  );
  mux_cell mux94 (
    .a (net161),
    .b (net159),
    .sel (net23),
    .out (net163)
  );
  mux_cell mux95 (
    .a (net161),
    .b (net159),
    .sel (net23),
    .out (net164)
  );
  mux_cell mux96 (
    .a (net160),
    .b (net162),
    .sel (net25),
    .out (net165)
  );
  mux_cell mux97 (
    .a (net163),
    .b (net164),
    .sel (net25),
    .out (net166)
  );
  mux_cell mux98 (
    .a (net165),
    .b (net166),
    .sel (net27),
    .out (net167)
  );
  mux_cell mux99 (
    .a (net168),
    .b (net168),
    .sel (net23),
    .out (net169)
  );
  mux_cell mux100 (
    .a (net168),
    .b (net168),
    .sel (net23),
    .out (net170)
  );
  mux_cell mux101 (
    .a (net168),
    .b (net168),
    .sel (net23),
    .out (net171)
  );
  mux_cell mux102 (
    .a (net172),
    .b (net172),
    .sel (net23),
    .out (net173)
  );
  mux_cell mux103 (
    .a (net169),
    .b (net170),
    .sel (net25),
    .out (net174)
  );
  mux_cell mux104 (
    .a (net171),
    .b (net173),
    .sel (net25),
    .out (net175)
  );
  mux_cell mux105 (
    .a (net174),
    .b (net175),
    .sel (net27),
    .out (net176)
  );
  mux_cell mux106 (
    .a (net177),
    .b (net177),
    .sel (net23),
    .out (net178)
  );
  mux_cell mux107 (
    .a (net179),
    .b (net179),
    .sel (net23),
    .out (net180)
  );
  mux_cell mux108 (
    .a (net177),
    .b (net177),
    .sel (net23),
    .out (net181)
  );
  mux_cell mux109 (
    .a (net177),
    .b (net179),
    .sel (net23),
    .out (net182)
  );
  mux_cell mux110 (
    .a (net178),
    .b (net180),
    .sel (net25),
    .out (net183)
  );
  mux_cell mux111 (
    .a (net181),
    .b (net182),
    .sel (net25),
    .out (net184)
  );
  mux_cell mux112 (
    .a (net183),
    .b (net184),
    .sel (net27),
    .out (net185)
  );
  mux_cell mux113 (
    .a (net186),
    .b (net186),
    .sel (net23),
    .out (net187)
  );
  mux_cell mux114 (
    .a (net186),
    .b (net188),
    .sel (net23),
    .out (net189)
  );
  mux_cell mux115 (
    .a (net188),
    .b (net186),
    .sel (net23),
    .out (net190)
  );
  mux_cell mux116 (
    .a (net186),
    .b (net188),
    .sel (net23),
    .out (net191)
  );
  mux_cell mux117 (
    .a (net187),
    .b (net189),
    .sel (net25),
    .out (net192)
  );
  mux_cell mux118 (
    .a (net190),
    .b (net191),
    .sel (net25),
    .out (net193)
  );
  mux_cell mux119 (
    .a (net192),
    .b (net193),
    .sel (net27),
    .out (net194)
  );
  mux_cell mux120 (
    .a (net195),
    .b (net195),
    .sel (net23),
    .out (net196)
  );
  mux_cell mux121 (
    .a (net195),
    .b (net195),
    .sel (net23),
    .out (net197)
  );
  mux_cell mux122 (
    .a (net198),
    .b (net195),
    .sel (net23),
    .out (net199)
  );
  mux_cell mux123 (
    .a (net198),
    .b (net195),
    .sel (net23),
    .out (net200)
  );
  mux_cell mux124 (
    .a (net196),
    .b (net197),
    .sel (net25),
    .out (net201)
  );
  mux_cell mux125 (
    .a (net199),
    .b (net200),
    .sel (net25),
    .out (net202)
  );
  mux_cell mux126 (
    .a (net201),
    .b (net202),
    .sel (net27),
    .out (net203)
  );
  mux_cell mux127 (
    .a (net204),
    .b (net205),
    .sel (net23),
    .out (net206)
  );
  mux_cell mux128 (
    .a (net204),
    .b (net204),
    .sel (net23),
    .out (net207)
  );
  mux_cell mux129 (
    .a (net205),
    .b (net204),
    .sel (net23),
    .out (net208)
  );
  mux_cell mux130 (
    .a (net204),
    .b (net205),
    .sel (net23),
    .out (net209)
  );
  mux_cell mux131 (
    .a (net206),
    .b (net207),
    .sel (net25),
    .out (net210)
  );
  mux_cell mux132 (
    .a (net208),
    .b (net209),
    .sel (net25),
    .out (net211)
  );
  mux_cell mux133 (
    .a (net210),
    .b (net211),
    .sel (net27),
    .out (net212)
  );
  mux_cell mux134 (
    .a (net213),
    .b (net213),
    .sel (net23),
    .out (net214)
  );
  mux_cell mux135 (
    .a (net213),
    .b (net215),
    .sel (net23),
    .out (net216)
  );
  mux_cell mux136 (
    .a (net215),
    .b (net215),
    .sel (net23),
    .out (net217)
  );
  mux_cell mux137 (
    .a (net215),
    .b (net213),
    .sel (net23),
    .out (net218)
  );
  mux_cell mux138 (
    .a (net214),
    .b (net216),
    .sel (net25),
    .out (net219)
  );
  mux_cell mux139 (
    .a (net217),
    .b (net218),
    .sel (net25),
    .out (net220)
  );
  mux_cell mux140 (
    .a (net219),
    .b (net220),
    .sel (net27),
    .out (net221)
  );
  mux_cell mux141 (
    .a (net222),
    .b (net222),
    .sel (net23),
    .out (net223)
  );
  mux_cell mux142 (
    .a (net224),
    .b (net224),
    .sel (net23),
    .out (net225)
  );
  mux_cell mux143 (
    .a (net224),
    .b (net222),
    .sel (net23),
    .out (net226)
  );
  mux_cell mux144 (
    .a (net222),
    .b (net222),
    .sel (net23),
    .out (net227)
  );
  mux_cell mux145 (
    .a (net223),
    .b (net225),
    .sel (net25),
    .out (net228)
  );
  mux_cell mux146 (
    .a (net226),
    .b (net227),
    .sel (net25),
    .out (net229)
  );
  mux_cell mux147 (
    .a (net228),
    .b (net229),
    .sel (net27),
    .out (net230)
  );
  mux_cell mux148 (
    .a (net231),
    .b (net231),
    .sel (net23),
    .out (net232)
  );
  mux_cell mux149 (
    .a (net233),
    .b (net233),
    .sel (net23),
    .out (net234)
  );
  mux_cell mux150 (
    .a (net231),
    .b (net231),
    .sel (net23),
    .out (net235)
  );
  mux_cell mux151 (
    .a (net231),
    .b (net231),
    .sel (net23),
    .out (net236)
  );
  mux_cell mux152 (
    .a (net232),
    .b (net234),
    .sel (net25),
    .out (net237)
  );
  mux_cell mux153 (
    .a (net235),
    .b (net236),
    .sel (net25),
    .out (net238)
  );
  mux_cell mux154 (
    .a (net237),
    .b (net238),
    .sel (net27),
    .out (net239)
  );
  mux_cell mux155 (
    .a (net240),
    .b (net241),
    .sel (net23),
    .out (net242)
  );
  mux_cell mux156 (
    .a (net240),
    .b (net240),
    .sel (net23),
    .out (net243)
  );
  mux_cell mux157 (
    .a (net240),
    .b (net241),
    .sel (net23),
    .out (net244)
  );
  mux_cell mux158 (
    .a (net241),
    .b (net241),
    .sel (net23),
    .out (net245)
  );
  mux_cell mux159 (
    .a (net242),
    .b (net243),
    .sel (net25),
    .out (net246)
  );
  mux_cell mux160 (
    .a (net244),
    .b (net245),
    .sel (net25),
    .out (net247)
  );
  mux_cell mux161 (
    .a (net246),
    .b (net247),
    .sel (net27),
    .out (net248)
  );
  mux_cell mux162 (
    .a (net249),
    .b (net250),
    .sel (net23),
    .out (net251)
  );
  mux_cell mux163 (
    .a (net250),
    .b (net249),
    .sel (net23),
    .out (net252)
  );
  mux_cell mux164 (
    .a (net250),
    .b (net250),
    .sel (net23),
    .out (net253)
  );
  mux_cell mux165 (
    .a (net249),
    .b (net250),
    .sel (net23),
    .out (net254)
  );
  mux_cell mux166 (
    .a (net251),
    .b (net252),
    .sel (net25),
    .out (net255)
  );
  mux_cell mux168 (
    .a (net255),
    .b (net256),
    .sel (net27),
    .out (net257)
  );
  mux_cell mux169 (
    .a (net258),
    .b (net259),
    .sel (net23),
    .out (net260)
  );
  mux_cell mux170 (
    .a (net259),
    .b (net259),
    .sel (net23),
    .out (net261)
  );
  mux_cell mux171 (
    .a (net258),
    .b (net259),
    .sel (net23),
    .out (net262)
  );
  mux_cell mux172 (
    .a (net259),
    .b (net258),
    .sel (net23),
    .out (net263)
  );
  mux_cell mux173 (
    .a (net260),
    .b (net261),
    .sel (net25),
    .out (net264)
  );
  mux_cell mux174 (
    .a (net262),
    .b (net263),
    .sel (net25),
    .out (net265)
  );
  mux_cell mux175 (
    .a (net264),
    .b (net265),
    .sel (net27),
    .out (net266)
  );
  mux_cell mux176 (
    .a (net267),
    .b (net267),
    .sel (net23),
    .out (net268)
  );
  mux_cell mux177 (
    .a (net269),
    .b (net267),
    .sel (net23),
    .out (net270)
  );
  mux_cell mux178 (
    .a (net267),
    .b (net269),
    .sel (net23),
    .out (net271)
  );
  mux_cell mux179 (
    .a (net267),
    .b (net269),
    .sel (net23),
    .out (net272)
  );
  mux_cell mux180 (
    .a (net268),
    .b (net270),
    .sel (net25),
    .out (net273)
  );
  mux_cell mux181 (
    .a (net271),
    .b (net272),
    .sel (net25),
    .out (net274)
  );
  mux_cell mux182 (
    .a (net273),
    .b (net274),
    .sel (net27),
    .out (net275)
  );
  mux_cell mux183 (
    .a (net276),
    .b (net276),
    .sel (net23),
    .out (net277)
  );
  mux_cell mux184 (
    .a (net276),
    .b (net276),
    .sel (net23),
    .out (net278)
  );
  mux_cell mux185 (
    .a (net276),
    .b (net276),
    .sel (net23),
    .out (net279)
  );
  mux_cell mux186 (
    .a (net276),
    .b (net276),
    .sel (net23),
    .out (net280)
  );
  mux_cell mux187 (
    .a (net277),
    .b (net278),
    .sel (net25),
    .out (net281)
  );
  mux_cell mux188 (
    .a (net279),
    .b (net280),
    .sel (net25),
    .out (net282)
  );
  mux_cell mux189 (
    .a (net281),
    .b (net282),
    .sel (net27),
    .out (net283)
  );
  mux_cell mux190 (
    .a (net284),
    .b (net284),
    .sel (net23),
    .out (net285)
  );
  mux_cell mux191 (
    .a (net284),
    .b (net286),
    .sel (net23),
    .out (net287)
  );
  mux_cell mux192 (
    .a (net284),
    .b (net284),
    .sel (net23),
    .out (net288)
  );
  mux_cell mux193 (
    .a (net284),
    .b (net284),
    .sel (net23),
    .out (net289)
  );
  mux_cell mux194 (
    .a (net285),
    .b (net287),
    .sel (net25),
    .out (net290)
  );
  mux_cell mux195 (
    .a (net288),
    .b (net289),
    .sel (net25),
    .out (net291)
  );
  mux_cell mux196 (
    .a (net290),
    .b (net291),
    .sel (net27),
    .out (net292)
  );
  mux_cell mux197 (
    .a (net293),
    .b (net293),
    .sel (net23),
    .out (net294)
  );
  mux_cell mux198 (
    .a (net293),
    .b (net293),
    .sel (net23),
    .out (net295)
  );
  mux_cell mux199 (
    .a (net293),
    .b (net293),
    .sel (net23),
    .out (net296)
  );
  mux_cell mux200 (
    .a (net297),
    .b (net293),
    .sel (net23),
    .out (net298)
  );
  mux_cell mux201 (
    .a (net294),
    .b (net295),
    .sel (net25),
    .out (net299)
  );
  mux_cell mux202 (
    .a (net296),
    .b (net298),
    .sel (net25),
    .out (net300)
  );
  mux_cell mux203 (
    .a (net299),
    .b (net300),
    .sel (net27),
    .out (net301)
  );
  mux_cell mux204 (
    .a (net302),
    .b (net302),
    .sel (net23),
    .out (net303)
  );
  mux_cell mux205 (
    .a (net302),
    .b (net302),
    .sel (net23),
    .out (net304)
  );
  mux_cell mux206 (
    .a (net302),
    .b (net302),
    .sel (net23),
    .out (net305)
  );
  mux_cell mux207 (
    .a (net302),
    .b (net306),
    .sel (net23),
    .out (net307)
  );
  mux_cell mux208 (
    .a (net303),
    .b (net304),
    .sel (net25),
    .out (net308)
  );
  mux_cell mux209 (
    .a (net305),
    .b (net307),
    .sel (net25),
    .out (net309)
  );
  mux_cell mux210 (
    .a (net308),
    .b (net309),
    .sel (net27),
    .out (net310)
  );
  mux_cell mux211 (
    .a (net311),
    .b (net312),
    .sel (net23),
    .out (net313)
  );
  mux_cell mux212 (
    .a (net312),
    .b (net311),
    .sel (net23),
    .out (net314)
  );
  mux_cell mux213 (
    .a (net311),
    .b (net311),
    .sel (net23),
    .out (net315)
  );
  mux_cell mux214 (
    .a (net311),
    .b (net312),
    .sel (net23),
    .out (net316)
  );
  mux_cell mux215 (
    .a (net313),
    .b (net314),
    .sel (net25),
    .out (net317)
  );
  mux_cell mux216 (
    .a (net315),
    .b (net316),
    .sel (net25),
    .out (net318)
  );
  mux_cell mux217 (
    .a (net317),
    .b (net318),
    .sel (net27),
    .out (net319)
  );
  mux_cell mux218 (
    .a (net320),
    .b (net321),
    .sel (net23),
    .out (net322)
  );
  mux_cell mux219 (
    .a (net320),
    .b (net320),
    .sel (net23),
    .out (net323)
  );
  mux_cell mux220 (
    .a (net320),
    .b (net321),
    .sel (net23),
    .out (net324)
  );
  mux_cell mux221 (
    .a (net320),
    .b (net320),
    .sel (net23),
    .out (net325)
  );
  mux_cell mux222 (
    .a (net322),
    .b (net323),
    .sel (net25),
    .out (net326)
  );
  mux_cell mux223 (
    .a (net324),
    .b (net325),
    .sel (net25),
    .out (net327)
  );
  mux_cell mux224 (
    .a (net326),
    .b (net327),
    .sel (net27),
    .out (net328)
  );
  mux_cell mux167 (
    .a (net50),
    .b (net59),
    .sel (net3),
    .out (net329)
  );
  mux_cell mux225 (
    .a (net68),
    .b (net77),
    .sel (net3),
    .out (net330)
  );
  mux_cell mux226 (
    .a (net86),
    .b (net95),
    .sel (net3),
    .out (net331)
  );
  mux_cell mux227 (
    .a (net104),
    .b (net113),
    .sel (net3),
    .out (net332)
  );
  mux_cell mux228 (
    .a (net329),
    .b (net330),
    .sel (net4),
    .out (net333)
  );
  mux_cell mux229 (
    .a (net331),
    .b (net332),
    .sel (net4),
    .out (net334)
  );
  mux_cell mux230 (
    .a (net333),
    .b (net334),
    .sel (net5),
    .out (net335)
  );
  mux_cell mux231 (
    .a (net122),
    .b (net131),
    .sel (net3),
    .out (net336)
  );
  mux_cell mux232 (
    .a (net140),
    .b (net149),
    .sel (net3),
    .out (net337)
  );
  mux_cell mux233 (
    .a (net158),
    .b (net167),
    .sel (net3),
    .out (net338)
  );
  mux_cell mux234 (
    .a (net176),
    .b (net185),
    .sel (net3),
    .out (net339)
  );
  mux_cell mux235 (
    .a (net336),
    .b (net337),
    .sel (net4),
    .out (net340)
  );
  mux_cell mux236 (
    .a (net338),
    .b (net339),
    .sel (net4),
    .out (net341)
  );
  mux_cell mux237 (
    .a (net340),
    .b (net341),
    .sel (net5),
    .out (net342)
  );
  mux_cell mux238 (
    .a (net194),
    .b (net203),
    .sel (net3),
    .out (net343)
  );
  mux_cell mux239 (
    .a (net212),
    .b (net221),
    .sel (net3),
    .out (net344)
  );
  mux_cell mux240 (
    .a (net230),
    .b (net239),
    .sel (net3),
    .out (net345)
  );
  mux_cell mux241 (
    .a (net248),
    .b (net257),
    .sel (net3),
    .out (net346)
  );
  mux_cell mux242 (
    .a (net343),
    .b (net344),
    .sel (net4),
    .out (net347)
  );
  mux_cell mux243 (
    .a (net345),
    .b (net346),
    .sel (net4),
    .out (net348)
  );
  mux_cell mux244 (
    .a (net347),
    .b (net348),
    .sel (net5),
    .out (net349)
  );
  mux_cell mux245 (
    .a (net266),
    .b (net275),
    .sel (net3),
    .out (net350)
  );
  mux_cell mux246 (
    .a (net283),
    .b (net292),
    .sel (net3),
    .out (net351)
  );
  mux_cell mux247 (
    .a (net301),
    .b (net310),
    .sel (net3),
    .out (net352)
  );
  mux_cell mux248 (
    .a (net319),
    .b (net328),
    .sel (net3),
    .out (net353)
  );
  mux_cell mux249 (
    .a (net350),
    .b (net351),
    .sel (net4),
    .out (net354)
  );
  mux_cell mux250 (
    .a (net352),
    .b (net353),
    .sel (net4),
    .out (net355)
  );
  mux_cell mux251 (
    .a (net354),
    .b (net355),
    .sel (net5),
    .out (net356)
  );
  mux_cell mux256 (
    .a (net335),
    .b (net342),
    .sel (net6),
    .out (net357)
  );
  mux_cell mux257 (
    .a (net349),
    .b (net356),
    .sel (net6),
    .out (net358)
  );
  mux_cell mux258 (
    .a (net357),
    .b (net358),
    .sel (net7),
    .out (net41)
  );
  mux_cell mux252 (
    .a (net253),
    .b (net254),
    .sel (net25),
    .out (net256)
  );
endmodule
